`timescale 1ps/1ps

`include "../data_macros.sv"

module generate_ray (
    input wire clk,
    input wire rst_n,
    input 

);
    
endmodule
