`ifndef DATA_MACROS_SV
`define DATA_MACROS_SV

`define LAMBERTIAN 2'd0
`define MIRROR     2'd1

`define INFINITY_24             24'h7FFFFF
`define NEGATIVE_INFINITY_24    24'h800000

`endif
